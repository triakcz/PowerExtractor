SPEED SENSE

.SUBCKT BCV47 1 2 3
*
* For use with Microsim PSPICE 
* please modify the AREA statement
* in this model:  e.g.
* SPICE: 
* Q2 1 22 3 BCV27 AREA = 5.1 
* PSPICE:
* Q2 1 22 3 BCV27 5.1 
* VTF, ITF, XTF are set to 
* default values 
*
Q1 1 2 33 BCV47 1 
Q2 1 33 3 BCV47 5.1 
.ENDS BCV47

*
.MODEL BCV47 NPN 
+ IS = 1.35E-14 
+ NF = 0.9889 
+ ISE = 4.441E-28 
+ NE = 1.03 
+ BF = 204 
+ IKF = 0.1 
+ VAF = 94 
+ NR = 1 
+ ISC = 1E-32 
+ NC = 2 
+ BR = 5 
+ IKR = 0.1 
+ VAR = 10 
+ RB = 45 
+ IRB = 7E-06 
+ RBM = 1 
+ RE = 0.25 
+ RC = 2 
+ XTB = 0 
+ EG = 1.11 
+ XTI = 3 
+ CJE = 1.445E-11 
+ VJE = 0.9 
+ MJE = 0.3635 
+ TF = 7E-10 
+ XTF = 1 
+ VTF = 1000 
+ ITF = 0.01 
+ PTF = 0 
+ CJC = 4.89E-12 
+ VJC = 0.6559 
+ MJC = 0.5115 
+ XCJC = 1 
+ TR = 1E-07 
+ CJS = 0 
+ VJS = 0.75 
+ MJS = 0.333 
+ FC = 0.999

.MODEL 1N4148 D 
+ IS = 4.352E-9 
+ N = 1.906 
+ BV = 110 
+ IBV = 0.0001 
+ RS = 0.6458 
+ CJO = 7.048E-13 
+ VJ = 0.869 
+ M = 0.03 
+ FC = 0.5 
+ TT = 3.48E-9 

Vdyn	1	2	SIN (	0	10	80	0	0	0)
V5	9	0	DC	5V
D1	0	1	1N4148
D2	0	2	1N4148
D5	1	3	1N4148
D6	2	4	1N4148
R4	3	6	100k
R3	4	5	100k
R1	6	0	100k
R2	5	0	100k
R5	9	7	10k
R6	9	8	10k
R7	7	5	100k
R8	8	6	100k
X1	7	6	0	BCV47
X2	8	5	0	BCV47



